VERSION 5.6 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 2000 ;
END UNITS

MANUFACTURINGGRID 0.000500 ; 

CLEARANCEMEASURE EUCLIDEAN ; 

USEMINSPACING OBS ON ; 

SITE CoreSite
    CLASS CORE ;
    SIZE 2.400000 BY 2.400000 ;
END CoreSite

LAYER m1
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 1.200000 ;
   AREA 0.810000 ;
   WIDTH 1.200000 ;
   SPACING 1.200000 ;
   PITCH 2.400000 2.400000 ;
END m1

LAYER v1
    TYPE CUT ;
    SPACING 0.900000 ;
    WIDTH 0.600000 ;
END v1

LAYER m2
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 1.200000 ;
   AREA 0.810000 ;
   WIDTH 1.200000 ;
   SPACING 1.200000 ;
   PITCH 2.400000 2.400000 ;
END m2

LAYER v2
    TYPE CUT ;
    SPACING 0.900000 ;
    WIDTH 0.600000 ;
END v2

LAYER m3
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 1.800000 ;
   AREA 2.250000 ;
   WIDTH 1.800000 ;
   SPACING 1.200000 ;
   PITCH 3.000000 3.000000 ;
END m3

LAYER v3
    TYPE CUT ;
    SPACING 0.900000 ;
    WIDTH 0.600000 ;
END v3

LAYER m4
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 1.200000 ;
   AREA 0.810000 ;
   WIDTH 1.200000 ;
   SPACING 1.200000 ;
   PITCH 2.400000 2.400000 ;
END m4

LAYER v4
    TYPE CUT ;
    SPACING 0.900000 ;
    WIDTH 0.600000 ;
END v4

LAYER m5
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 1.800000 ;
   AREA 2.250000 ;
   WIDTH 1.800000 ;
   SPACING 1.200000 ;
   PITCH 3.000000 3.000000 ;
END m5


VIA v1_C DEFAULT
   LAYER m1 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER v1 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
   LAYER m2 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
END v1_C

VIA v2_C DEFAULT
   LAYER m2 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER v2 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
   LAYER m3 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
END v2_C

VIA v3_C DEFAULT
   LAYER m3 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER v3 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
   LAYER m4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
END v3_C

VIA v4_C DEFAULT
   LAYER m4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER v4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
   LAYER m5 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
END v4_C

MACRO _0_0cell_0_0g1x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g1x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 7.200000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g1x0

MACRO _0_0cell_0_0g1x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g1x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 7.200000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g1x0_plug

MACRO _0_0cell_0_0g0x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 28.800000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 14.400000 6.000000 15.600000 7.200000 ;
        END
    END in_51_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g0x0

MACRO _0_0cell_0_0g0x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 28.800000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 14.400000 6.000000 15.600000 7.200000 ;
        END
    END in_51_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g0x0_plug

MACRO _0_0cell_0_0g2x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g2x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 48.000000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 9.600000 6.000000 10.800000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 16.800000 6.000000 18.000000 7.200000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 24.000000 6.000000 25.200000 7.200000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 31.200000 6.000000 32.400000 7.200000 ;
        END
    END in_54_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g2x0

MACRO _0_0cell_0_0g2x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g2x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 48.000000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 9.600000 6.000000 10.800000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 16.800000 6.000000 18.000000 7.200000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 24.000000 6.000000 25.200000 7.200000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 31.200000 6.000000 32.400000 7.200000 ;
        END
    END in_54_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g2x0_plug

MACRO _0_0cell_0_0g5x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g5x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 12.000000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 4.800000 6.000000 6.000000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 7.200000 6.000000 8.400000 7.200000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g5x0

MACRO _0_0cell_0_0g5x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g5x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 12.000000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 4.800000 6.000000 6.000000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 7.200000 6.000000 8.400000 7.200000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g5x0_plug

MACRO _0_0cell_0_0g3x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g3x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 60.000000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 12.000000 6.000000 13.200000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 21.600000 6.000000 22.800000 7.200000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 31.200000 6.000000 32.400000 7.200000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 40.800000 6.000000 42.000000 7.200000 ;
        END
    END in_54_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g3x0

MACRO _0_0cell_0_0g3x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g3x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 60.000000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 12.000000 6.000000 13.200000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 21.600000 6.000000 22.800000 7.200000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 31.200000 6.000000 32.400000 7.200000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 40.800000 6.000000 42.000000 7.200000 ;
        END
    END in_54_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g3x0_plug

MACRO _0_0cell_0_0g4x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g4x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 72.000000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 14.400000 6.000000 15.600000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 26.400000 6.000000 27.600000 7.200000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 38.400000 6.000000 39.600000 7.200000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 50.400000 6.000000 51.600000 7.200000 ;
        END
    END in_54_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g4x0

MACRO _0_0cell_0_0g4x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g4x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 72.000000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 14.400000 6.000000 15.600000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 26.400000 6.000000 27.600000 7.200000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 38.400000 6.000000 39.600000 7.200000 ;
        END
    END in_53_6
    PIN in_54_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 50.400000 6.000000 51.600000 7.200000 ;
        END
    END in_54_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g4x0_plug

MACRO _0_0cell_0_0g8x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g8x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 36.000000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 9.600000 6.000000 10.800000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 16.800000 6.000000 18.000000 7.200000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 24.000000 6.000000 25.200000 7.200000 ;
        END
    END in_53_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g8x0

MACRO _0_0cell_0_0g8x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g8x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 36.000000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 9.600000 6.000000 10.800000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 16.800000 6.000000 18.000000 7.200000 ;
        END
    END in_52_6
    PIN in_53_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 24.000000 6.000000 25.200000 7.200000 ;
        END
    END in_53_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g8x0_plug

MACRO _0_0cell_0_0g6x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g6x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 31.200000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 9.600000 6.000000 10.800000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 16.800000 6.000000 18.000000 7.200000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g6x0

MACRO _0_0cell_0_0g6x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g6x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 31.200000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 9.600000 6.000000 10.800000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 16.800000 6.000000 18.000000 7.200000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g6x0_plug

MACRO _0_0cell_0_0g7x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g7x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 9.600000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 4.800000 6.000000 6.000000 7.200000 ;
        END
    END in_51_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g7x0

MACRO _0_0cell_0_0g7x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g7x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 9.600000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 4.800000 6.000000 6.000000 7.200000 ;
        END
    END in_51_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g7x0_plug

MACRO _0_0cell_0_0g9x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g9x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 28.800000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 9.600000 6.000000 10.800000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 16.800000 6.000000 18.000000 7.200000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g9x0

MACRO _0_0cell_0_0g9x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g9x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 28.800000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 9.600000 6.000000 10.800000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 16.800000 6.000000 18.000000 7.200000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g9x0_plug

MACRO _0_0cell_0_0g10x0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g10x0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 12.000000 BY 12.000000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 4.800000 6.000000 6.000000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 7.200000 6.000000 8.400000 7.200000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g10x0

MACRO _0_0cell_0_0g10x0_plug
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g10x0_plug 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 12.000000 BY 21.600000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 6.000000 3.600000 7.200000 ;
        END
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 4.800000 6.000000 6.000000 7.200000 ;
        END
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 7.200000 6.000000 8.400000 7.200000 ;
        END
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m2 ;
        RECT 2.400000 2.400000 3.600000 3.600000 ;
        END
    END out
END _0_0cell_0_0g10x0_plug

